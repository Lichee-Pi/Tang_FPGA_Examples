// Verilog netlist created by TD v4.2.217
// Wed Jul 25 16:58:49 2018

`timescale 1ns / 1ps
module img  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_rom.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [13:0] addra;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_rom.v(18)
  input clka;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_rom.v(19)
  input rsta;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_rom.v(20)
  output [15:0] doa;  // H:/Work/FPGA/AnLogic/LicheeTang/demo/test_lcd_camera/test_camera/project/al_ip/ip_rom.v(16)

  wire [0:2] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b0/B0_2 ;
  wire  \inst_doa_mux_b0/B0_3 ;
  wire  \inst_doa_mux_b0/B1_0 ;
  wire  \inst_doa_mux_b0/B1_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b1/B0_2 ;
  wire  \inst_doa_mux_b1/B0_3 ;
  wire  \inst_doa_mux_b1/B1_0 ;
  wire  \inst_doa_mux_b1/B1_1 ;
  wire  \inst_doa_mux_b10/B0_0 ;
  wire  \inst_doa_mux_b10/B0_1 ;
  wire  \inst_doa_mux_b10/B0_2 ;
  wire  \inst_doa_mux_b10/B0_3 ;
  wire  \inst_doa_mux_b10/B1_0 ;
  wire  \inst_doa_mux_b10/B1_1 ;
  wire  \inst_doa_mux_b11/B0_0 ;
  wire  \inst_doa_mux_b11/B0_1 ;
  wire  \inst_doa_mux_b11/B0_2 ;
  wire  \inst_doa_mux_b11/B0_3 ;
  wire  \inst_doa_mux_b11/B1_0 ;
  wire  \inst_doa_mux_b11/B1_1 ;
  wire  \inst_doa_mux_b12/B0_0 ;
  wire  \inst_doa_mux_b12/B0_1 ;
  wire  \inst_doa_mux_b12/B0_2 ;
  wire  \inst_doa_mux_b12/B0_3 ;
  wire  \inst_doa_mux_b12/B1_0 ;
  wire  \inst_doa_mux_b12/B1_1 ;
  wire  \inst_doa_mux_b13/B0_0 ;
  wire  \inst_doa_mux_b13/B0_1 ;
  wire  \inst_doa_mux_b13/B0_2 ;
  wire  \inst_doa_mux_b13/B0_3 ;
  wire  \inst_doa_mux_b13/B1_0 ;
  wire  \inst_doa_mux_b13/B1_1 ;
  wire  \inst_doa_mux_b14/B0_0 ;
  wire  \inst_doa_mux_b14/B0_1 ;
  wire  \inst_doa_mux_b14/B0_2 ;
  wire  \inst_doa_mux_b14/B0_3 ;
  wire  \inst_doa_mux_b14/B1_0 ;
  wire  \inst_doa_mux_b14/B1_1 ;
  wire  \inst_doa_mux_b15/B0_0 ;
  wire  \inst_doa_mux_b15/B0_1 ;
  wire  \inst_doa_mux_b15/B0_2 ;
  wire  \inst_doa_mux_b15/B0_3 ;
  wire  \inst_doa_mux_b15/B1_0 ;
  wire  \inst_doa_mux_b15/B1_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b2/B0_2 ;
  wire  \inst_doa_mux_b2/B0_3 ;
  wire  \inst_doa_mux_b2/B1_0 ;
  wire  \inst_doa_mux_b2/B1_1 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b3/B0_2 ;
  wire  \inst_doa_mux_b3/B0_3 ;
  wire  \inst_doa_mux_b3/B1_0 ;
  wire  \inst_doa_mux_b3/B1_1 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b4/B0_2 ;
  wire  \inst_doa_mux_b4/B0_3 ;
  wire  \inst_doa_mux_b4/B1_0 ;
  wire  \inst_doa_mux_b4/B1_1 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b5/B0_2 ;
  wire  \inst_doa_mux_b5/B0_3 ;
  wire  \inst_doa_mux_b5/B1_0 ;
  wire  \inst_doa_mux_b5/B1_1 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b6/B0_2 ;
  wire  \inst_doa_mux_b6/B0_3 ;
  wire  \inst_doa_mux_b6/B1_0 ;
  wire  \inst_doa_mux_b6/B1_1 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire  \inst_doa_mux_b7/B0_2 ;
  wire  \inst_doa_mux_b7/B0_3 ;
  wire  \inst_doa_mux_b7/B1_0 ;
  wire  \inst_doa_mux_b7/B1_1 ;
  wire  \inst_doa_mux_b8/B0_0 ;
  wire  \inst_doa_mux_b8/B0_1 ;
  wire  \inst_doa_mux_b8/B0_2 ;
  wire  \inst_doa_mux_b8/B0_3 ;
  wire  \inst_doa_mux_b8/B1_0 ;
  wire  \inst_doa_mux_b8/B1_1 ;
  wire  \inst_doa_mux_b9/B0_0 ;
  wire  \inst_doa_mux_b9/B0_1 ;
  wire  \inst_doa_mux_b9/B0_2 ;
  wire  \inst_doa_mux_b9/B0_3 ;
  wire  \inst_doa_mux_b9/B1_0 ;
  wire  \inst_doa_mux_b9/B1_1 ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i0_008;
  wire inst_doa_i0_009;
  wire inst_doa_i0_010;
  wire inst_doa_i0_011;
  wire inst_doa_i0_012;
  wire inst_doa_i0_013;
  wire inst_doa_i0_014;
  wire inst_doa_i0_015;
  wire inst_doa_i4_000;
  wire inst_doa_i4_001;
  wire inst_doa_i4_002;
  wire inst_doa_i4_003;
  wire inst_doa_i4_004;
  wire inst_doa_i4_005;
  wire inst_doa_i4_006;
  wire inst_doa_i4_007;
  wire inst_doa_i4_008;
  wire inst_doa_i4_009;
  wire inst_doa_i4_010;
  wire inst_doa_i4_011;
  wire inst_doa_i4_012;
  wire inst_doa_i4_013;
  wire inst_doa_i4_014;
  wire inst_doa_i4_015;

  reg_sr_as_w1 addra_pipe_b0 (
    .clk(clka),
    .d(addra[11]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[0]));
  reg_sr_as_w1 addra_pipe_b1 (
    .clk(clka),
    .d(addra[12]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[1]));
  reg_sr_as_w1 addra_pipe_b2 (
    .clk(clka),
    .d(addra[13]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[2]));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h033FFFFFFFFFFFFFFFE00001FC0FFFFFFFFFFFFFFFFF45041FFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFF0001F800381FFFFFFFFFFFFFF0001F00030FFFFFFFFFFFFFFF8000700),
    .INIT_02(256'hFC007C007FFFFFFFFFFE0000FF8007C00FFFFFFFFFFFF80003F800780FFFFFFF),
    .INIT_03(256'hFFFFFFFF81007FFC01FE00FFFFFFFFFFFC0001FFC01FE006FFFFFFFFFFC8000F),
    .INIT_04(256'h3FFFE0FFF01FFFFFFFFFFF0021FFFE0FFF00FFFFFFFFFFF80807FFE03FF00FFF),
    .INIT_05(256'hFFF0FFFFFFC00F81FFFBFFF83FFFFFFFFFFC0061FFFF0FFF81FFFFFFFFFFF000),
    .INIT_06(256'hBBFF00007FFFE7FC06BFFFFF057B6001FBFFFC3FF80FFFFFF8017800FFBFFFC3),
    .INIT_07(256'hFF000197BFFFFFFBEF0001FFFFFC000D77FFFE3FFF300007FFFE7E00C77FFFF0),
    .INIT_08(256'hFFFDFEFC003FFFFF800003FFFFFFFFEFC001FFFFD80020FDFFFFFFFDF8001FFF),
    .INIT_09(256'hFFEFFE00403FD7FDFFFCFE007FFFFFE00003FEFFFFFFFFC003FFFFDC00607F9F),
    .INIT_0A(256'hFFBFEBFFBFF01FFFFFFF80803FEFFFBFFFFF00FFF7FBF01403FEFFFFFFDFE007),
    .INIT_0B(256'hC3FFFFEFFE2003FBFFBFFFBFF83FFFFFFFC3003F9FFCFFFBFF81FFBFFFF80003),
    .INIT_0C(256'h001F7FFFFFFFFFE7BFFFFFFFA002F7FF5FFFFFFC3FFFFEFFE0001F7DFBFFFBFF),
    .INIT_0D(256'h7FFD3FFFFFFFF5A01DFF7DDFFFFFE3FFFFFFFC2002DFCFF3FF7FFEF3FFFFFFE0),
    .INIT_0E(256'hC01FFFFFF7FF3FFF83DFFFFFFE43FD07FEFFEFEFFFDFFFFFDFFE1840FFFFDFFF),
    .INIT_0F(256'hFF7F027FDFFF7F80D7FE7003FFDFF00BF3FFFFFE007FF023FFFFDF907E3FFFFF),
    .INIT_10(256'hFE60083F07F03EFF8001FFF7FFFE0097F07F01EFF7000FFDFFF7D00DFFC7003E),
    .INIT_11(256'hFCF7FF003FFFFFDD00043807FFAFBBC003FFFFFFE00085C07FC7FBEC007FFFFF),
    .INIT_12(256'hFFC78000CB403FEFFBFE00FFFFFDF8000C0003FFFF7FE017FFFF3DA000C2003F),
    .INIT_13(256'h21C03FFFF03FFFFFEB7FFFFE043FC2FBFF03FFFFFE501809E181F83FFFF01FFF),
    .INIT_14(256'hF0E00407FFF07803803FDFF0FFFFD89CBFFFDE801803FFFF0FFFFE4F1FFFF1E0),
    .INIT_15(256'h01803FEBFF7FA2000024007FE07006F83FEFFAD00000401FFE03C04E03FFFF0F),
    .INIT_16(256'hF40000380003FC018077FBFFFF40000110002FC01C237FBFFFF80000010007FF),
    .INIT_17(256'h0300042FBEFFFBE0C000C400003800B8FFF7FFBE48000200000BC0088FFF7FF7),
    .INIT_18(256'hFFF80081C201000500001FFFFFFF840004001000400000FFFFFFFC4200280100),
    .INIT_19(256'h004023000BFFFFFFD000200000008230019FDFFFFF000008000002000001FFDF),
    .INIT_1A(256'hC7FFFC00030000100000400FFEBFFFD400140002200008009FFFFFFF00028080),
    .INIT_1B(256'h800F00000023FFFFFFFF153F000022000010FFFCFFFFE102F0B03280000003FF),
    .INIT_1C(256'h3FEFFFFFF1BFF1F03F80802407FF7FFFFF81FF0F80702000CDFFFFFFFFF0FFF0),
    .INIT_1D(256'hE31FC3FC0000181FDFFFFFF40FF1FE1FC02001C3FCFFFFFF831F1F01FC03F80C),
    .INIT_1E(256'hE3C02FFFFFFEEC3E3F04FE01F83C007FFFFFEF97F81F7FE06F81807BFFFFFFC0),
    .INIT_1F(256'h8FF181FFFEF97F3FC10BFFFFFCFE381FEF5F0FFCFC007FFFFFCFCFE3FFFFF07F),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n63,open_n64,addra[13]}),
    .dia({open_n68,open_n69,open_n70,open_n71,open_n72,open_n73,open_n74,1'b0,open_n75}),
    .rsta(rsta),
    .doa({open_n90,open_n91,open_n92,open_n93,open_n94,open_n95,open_n96,open_n97,inst_doa_i0_000}));
  // address_offset=0;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBAFBFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFF),
    .INIT_03(256'hFFFFFFFF80FFFFFFFFFFFF03FFFFFFFFFC3FFFFFFFFFFFF8FFFFFFFFFFC7FFFF),
    .INIT_04(256'hFFFFFFFFFFE001FFFFFFFF001FFFFFFFFFFF003FFFFFFFF007FFFFFFFFFFF00F),
    .INIT_05(256'h000C7FFFFFC004BFFFFFFFFFC0001FFFFFFC000BFFFFFFFFFE0007FFFFFFE000),
    .INIT_06(256'h8071FFFFFFFFF803F83FFFFF00871FFFFFFFFFC007C7FFFFF8021FFFFFFFFFFC),
    .INIT_07(256'hFFFFFE001FFFE003F0FFFFFFFFF1FFF803FFFE401F0FFFFFFFFF81FFC0FFFFF0),
    .INIT_08(256'hFC03FE03FFFFFFFFFFFE0007FFC00FE07FFFFFFFFFFFF081FFFC007F07FFFFFF),
    .INIT_09(256'hFFFFFFFFC0000FFC0FFD01FFFFFFFFFFFC0000FFC07FE03FFFFFFFFFFFE0001F),
    .INIT_0A(256'h007FC3FFC00FFFFFFFFFFF000013FC3FFC00FFFFFFFFFFEC00007FC1FFC01FFF),
    .INIT_0B(256'h3FFFFFFFFFC002003FFFFF8007FFFFFFFFFE000003F9FFF8007FFFFFFFFFE000),
    .INIT_0C(256'h000003FFFFF8001FFFFFFFFF6002001FDFFF8003FFFFFFFFFC000001FFFFF800),
    .INIT_0D(256'h0000FFFFFFFFFC200201FDFFF0001FFFFFFFFE0001000FF7FF0001FFFFFFFFF8),
    .INIT_0E(256'hEF80008007FFFF00001FFFFFFFB8008000FDFFE00003FFFFFFFF8040000FDFFF),
    .INIT_0F(256'hFF6200003FFFFFFF8001F007EFFE000007FFFFFDF80008207FFFE00000FFFFFF),
    .INIT_10(256'hFFFFF841FFF07FFF8002000FFFFFFF8007FE07EFFE000001FFFFFFF8803F007E),
    .INIT_11(256'hFDFFFE0080000FFF7FF807FFFF3FFBE0000001FFFFFF803FFFC5FBEC0000003F),
    .INIT_12(256'h001F7FFF81FFFFFDFFFE00000003FBFFF80FFFFFFF7FE00000007FDFFF80FFFF),
    .INIT_13(256'hFFFFFFFBF000000002C00000FFFFFFFBFF000000007FFFFA0EFDFFFFFFE02000),
    .INIT_14(256'h007FF880000F07FFFFFFFFF000001FFC0000A0FFFFFFFFFF0800000F4000060F),
    .INIT_15(256'hFC7FC01FFFFF83FFFFF780001F87F807BFEFFA00FFFFD80000F8BFB3FBFFFF00),
    .INIT_16(256'hF2FFFFF9F80103FF778007FFFF1FFFFF9F80003FE3D8807FFFFFFFFFFD780000),
    .INIT_17(256'h007FFBD001FFFFE73FFFC7F00007FF47400FFFFE37FFFE3F00007FF77000FFFF),
    .INIT_18(256'hFFF83FFF43FF0003FFFDE001FFFF87FFFC0FF0000FFFFE002FFFBC7DFFF87F00),
    .INIT_19(256'hE07FFEFFF4003FFFF03FFC07FE00FFDFFE4003FFFD03FFE03FE001FFFFFE001F),
    .INIT_1A(256'h0FFFFE03FFE1FFFFFFFFFFF0007FFFE03FE40FFE3FFFF7FF8007FFFE03FD80FF),
    .INIT_1B(256'h0000FFFFFFDFC03FFFFF06FFF8000FFFFFFF7802FFFFF33DFF3801FFFFFDFD80),
    .INIT_1C(256'h7E07FFFFF07FFE00007FFFC8FFC07FFFFF03FFF00007FFFF77FC07FFFFF04FFF),
    .INIT_1D(256'hFF800003FE001FEE3FFFFFFBFFFC00003FF000FFE1FFFFFF9DFFE00007FF100F),
    .INIT_1E(256'h03FFF7FFFFFFF3FF800001FC003FFF3FFFFFFF6FF800001FC003FFF3FFFFFFFE),
    .INIT_1F(256'hFFFFFE000107007BFFB3FFFFFFFDFFC00000F0007FFF7FFFFFFFB7FC00000FC0),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n123,open_n124,addra[13]}),
    .dia({open_n128,open_n129,open_n130,open_n131,open_n132,open_n133,open_n134,1'b0,open_n135}),
    .rsta(rsta),
    .doa({open_n150,open_n151,open_n152,open_n153,open_n154,open_n155,open_n156,open_n157,inst_doa_i0_001}));
  // address_offset=0;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'h7FFFFFFFFFFFFFFFFFFFFFFFFEFF7FFFFFFFFFFFFFFBFFFFFFFDFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFF7FFFFFFBFFFFFFFFFFFFFFFFFBFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFE3FFBFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFBFFFF7FFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFDFC3FFFFFFFFFFFFFFFFFFFFFFFC3FFFFFBFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFF03FFFFFFFFFFFFFFFFFF9FFDF01FDFFFFFFFFFFFFFFFFFFFFF83FBFFFFFF),
    .INIT_0D(256'hFFFDFFFFFFFFE01FFE00FDFFFFFFFFFFFFFFFF9FFEE01FF7FFFFFFFFFFFFFFFF),
    .INIT_0E(256'hF060000007FFFEFFC3FFFFFFFF84007800FFFFEFFF1FFFFFFFFC403FC00FDFFF),
    .INIT_0F(256'hFF7C00FFFFFFFFC070019FFFEFFFF807FFFFFFFC07000FE07FFFFFE07FFFFFFF),
    .INIT_10(256'hFFC007C1F80FFFFF8001FFFFFFFE00780781FBFFFD001FFFFFFFF0078038FFFE),
    .INIT_11(256'h01F700007FFFFFFF8007C7FC00FFF80007FFFFFFF8007C3F8039FBE0003FFFFF),
    .INIT_12(256'hFFFF0000787FC003F80001FFFFFFFC0007EFFC001FC0000FFFFFFFE0007EFFC0),
    .INIT_13(256'h1E003FF8007FFFFFFC3FFF8007C003FF0003FFFFFFE0000600FE003FE0101FFF),
    .INIT_14(256'hFFFFFF07FFF00800003FFF00FFFFFFF0FFFF00006003FFE007FFFFF79FFFF800),
    .INIT_15(256'h0001FFE7FFFF3BFFFFF800FFE0000FF87FEFE1FEFFFFA01FFF00003C07FFFC9F),
    .INIT_16(256'hF7FFFFF60001FC0007FFFFFFFF7FFFFFE0003FC0003FFFBFFFFBFFFFFE8007FE),
    .INIT_17(256'h018003FFFFFFFFE7FFFFB8000038003FBFFFFFFE7FFFFFC000078001FFFFFFFF),
    .INIT_18(256'hFFF83FFFBC0000000001FFFFFFFF87FFFFF0000000003FFFDFFFFC7FFFF78000),
    .INIT_19(256'h000000000FFFFFFFF03FFFF80000000001FFFFFFFF03FFF7C0000000001FFFDF),
    .INIT_1A(256'hFFFFFF03F81E000000000007FFFFFFE03FFBF00000000000FFFFFFFE03FFFF00),
    .INIT_1B(256'h00070000001FFFDFFFFF07C00000300000007FFEFFFFF13F00400200000201FF),
    .INIT_1C(256'h7FF7FFFFF0C000000F8000007FFFBFFFFF00000000F8000007FFFBFFFFF07000),
    .INIT_1D(256'h000003FC000007FFFFFFFFFFE000001FC000007FFFFFFFFF3E000001F8002007),
    .INIT_1E(256'h003FF7FFFFFFFF000007FE000003FFFFFFFFFFF000003FE000007FFFFFFFFFFF),
    .INIT_1F(256'hFFF8000001F800043FC3FFFFFFFF8000007F000003FE7FFFFFFFF800001FF040),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n183,open_n184,addra[13]}),
    .dia({open_n188,open_n189,open_n190,open_n191,open_n192,open_n193,open_n194,1'b0,open_n195}),
    .rsta(rsta),
    .doa({open_n210,open_n211,open_n212,open_n213,open_n214,open_n215,open_n216,open_n217,inst_doa_i0_002}));
  // address_offset=0;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFEFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'h800FFFFFFFFFFFFFFF1FFFFFFF00FFFFFFFFFFFFFFF3FFFFFFFE07FFFFFFFFFF),
    .INIT_07(256'hFFFFFFF03FFFE0000FFFFFFFFFFFFFFF07FFFFC000FFFFFFFFFFFFFFF0FFFFFF),
    .INIT_08(256'hFC0001FFFFFFFFFFFFFFF807FFC0001FFFFFFFFFFFFFEF80FFFC0000FFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFC007FC0003FFFFFFFFFFFFFFF801FFC0001FFFFFFFFFFFFFFF803F),
    .INIT_0A(256'h01FFC4003FFFFFFFFFFFFFFFC00FFC0003FFFFFFFFFFFFFFFC00FFC0003FFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFE03FF80007FFFFFFFFFFFFFFFC03FFC0007FFFFFFFFFFFFFFFC),
    .INIT_0C(256'hFFE0FDFF0007FFFFFFFFFFFFFFFE0FFFC0007FFFFFFFFFFFFFFFE07DF80007FF),
    .INIT_0D(256'hFFFFFFFFFFFFE3FFF1FFFDC00FFFFFFFFFFFFF7FFF1FFFF000FFFFFFFFFFFFFF),
    .INIT_0E(256'hF01FFF7FFFFF81FFFFFFFFFFFF81FFF7FFFFF01FFFFFFFFFFFFC3FFF3FFFDE00),
    .INIT_0F(256'hFF9FFFFFFFFFFF800FFE6007EFE1FFFFFFFFFFFE00FFF41FFFFC1FFFFFFFFFFF),
    .INIT_10(256'hFFC0003E07F83FFFBFFFFFFFFFFE0007F87E07FFFBFFFFFFFFFFF0007FC7807E),
    .INIT_11(256'hFFF701FFFFFFFFFF00003803FF1FF81FFFFFFFFFF80003C07FE3FBE3FFFFFFFF),
    .INIT_12(256'hFFFF800001803FFFF801FFFFFFFFFC00001003FFFFC01FFFFFFFFFE00001003F),
    .INIT_13(256'hE1FFFFF80FFFFFFFFC000000F83FFFFF00FFFFFFFFE000000F03FFFFE00FFFFF),
    .INIT_14(256'hFF80000000000FFFFFFFFF0FFFFFE010000000FF9FFFFFE0FFFFFFF80000000F),
    .INIT_15(256'h007E001FFFFF7C00001000000007F007FFEFE7FF000000000000FFC3FFFFFC7F),
    .INIT_16(256'hF600001000000000780007FFFF4000000000000007C0007FFFF8000000000000),
    .INIT_17(256'h0000000000FFFFE78000000000000040000FFFFE700000000000000600007FFF),
    .INIT_18(256'hFFF83F000000000000000001FFFF87E000000000000000001FFFFC7C00100000),
    .INIT_19(256'h0000000000003FFFF03FC00000000000000003FFFF03F810000000000000003F),
    .INIT_1A(256'h0FFFFE03FC00000000000000007FFFE03FE00000000000000007FFFF03FE0000),
    .INIT_1B(256'h000000000000001FFFFF07C00000000000000001FFFFF13F0000000000000000),
    .INIT_1C(256'h800FFFFFF0C000000000000F80007FFFFF00000000000000000003FFFFF07000),
    .INIT_1D(256'h0000000001FFE0001FFFFFFFE0000000001FFF0000FFFFFF3E00000000001FF0),
    .INIT_1E(256'hFC000FFFFFFFFF0000000003FFC0007FFFFFFFF0000000003FFE0003FFFFFFFF),
    .INIT_1F(256'hFFF800000000FFC0000FFFFFFFFF8000000007FF8000FFFFFFFFF8000000003F),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n243,open_n244,addra[13]}),
    .dia({open_n248,open_n249,open_n250,open_n251,open_n252,open_n253,open_n254,1'b0,open_n255}),
    .rsta(rsta),
    .doa({open_n270,open_n271,open_n272,open_n273,open_n274,open_n275,open_n276,open_n277,inst_doa_i0_003}));
  // address_offset=0;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFF001FFFFFFFFFFFFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFFFF80FFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFE0007FFFFFFFFFFFFFFFFFFFFF000FFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFF800007FFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFC0003F),
    .INIT_0A(256'h003FFFFFFFFFFFFFFFFFFF000007FFFFFFFFFFFFFFFFFFF800007FFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFE000003FFFFFFFFFFFFFFFFFFE000003FFFFFFFFFFFFFFFFFFF000),
    .INIT_0C(256'h000001FCFFFFFFFFFFFFFFFFC000001FFFFFFFFFFFFFFFFFFC000003FFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFE0000000FE3FFFFFFFFFFFFFFF0000001FCFFFFFFFFFFFFFFFF8),
    .INIT_0E(256'hF00000000FE07FFFFFFFFFFFFF80000000FE0FFFFFFFFFFFFFFC0000000FE1FF),
    .INIT_0F(256'h00FFFFFFFFFFFF8000000007F01FFFFFFFFFFFFE000000007E03FFFFFFFFFFFF),
    .INIT_10(256'hFFC0000000003F007FFFFFFFFFFE0000000007F007FFFFFFFFFFF0000000007F),
    .INIT_11(256'h03F8FFFFFFFFFFFF00000000003F07FFFFFFFFFFF80000000003F41FFFFFFFFF),
    .INIT_12(256'hFFFF800000000003FFFFFFFFFFFFFC00000000003FBFFFFFFFFFFFE000000000),
    .INIT_13(256'h00003FC7FFFFFFFFFC000000000003FCFFFFFFFFFFE000000000003F9FFFFFFF),
    .INIT_14(256'hFFFFFC0000000000003FE0FFFFFFFFE0000000000003FC1FFFFFFFFF80000000),
    .INIT_15(256'h00000003FF00FFFFFFE00000000000003FF01FFFFFFF80000000000003FE03FF),
    .INIT_16(256'h09FFFFE000000000000007FF00BFFFFF800000000000007FF007FFFFFC000000),
    .INIT_17(256'h0000000000FFF8187FFF800000000000000FFF818FFFFC000000000000007FF8),
    .INIT_18(256'hFFC7C0FF8000000000000001FFFC781FFC000000000000001FFFC383FFE00000),
    .INIT_19(256'h0000000000003FFFEFC03C0000000000000003FFFEFC07E0000000000000003F),
    .INIT_1A(256'h0FFFFE3C0000000000000000007FFFE7C0000000000000000007FFFEFC018000),
    .INIT_1B(256'h000000000000001FFFFF08000000000000000000FFFFF0C00000000000000000),
    .INIT_1C(256'h000FFFFFF00000000000000000007FFFFF00000000000000000003FFFFF00000),
    .INIT_1D(256'h00000000000000001FFFFFF8000000000000000000FFFFFF0000000000000000),
    .INIT_1E(256'h00000FFFFFFFF000000000000000007FFFFFFE000000000000000003FFFFFFC0),
    .INIT_1F(256'hFFE00000000000000003FFFFFFFC00000000000000007FFFFFFF800000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n303,open_n304,addra[13]}),
    .dia({open_n308,open_n309,open_n310,open_n311,open_n312,open_n313,open_n314,1'b0,open_n315}),
    .rsta(rsta),
    .doa({open_n330,open_n331,open_n332,open_n333,open_n334,open_n335,open_n336,open_n337,inst_doa_i0_004}));
  // address_offset=0;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFDFFFFFFFFFFFFFFFEFFFEFFFFFFFFFFFFFFFFFFFFF36EFBBFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFC07FC0FFFFBFFFFFFFFFFFFFFF07FF0FFFF77FFFFFFFFFFFFFF87FF9FF),
    .INIT_02(256'h03FFFFFFFFFFFFFFFFFF007F807FFFFFFFFFFFFFFFFFF407FC07FFFBFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFC07C003FFFFFF77FFFFFFFFFFC07E003FFFFFF9FFFFFFFFFFF407F0),
    .INIT_04(256'h40001FFFF7FFFEFFFFFFFF7FE60003FFFE7FFFFFFFFFFFFFF078001FFFEFFFEF),
    .INIT_05(256'hFFE67FFFFFFFD03F000FFFFFFFFFFFFFFFFFFFF60000FFFFFDFFF7FFFFFFEFFE),
    .INIT_06(256'hC083FFFFBFFFDBFDFDBFFFFF3C405FFFC7FFFFFFFFF9FFFFFBFFC1FF00FFFFFF),
    .INIT_07(256'h00FFFE887FFFC00010FFFF0003FDFFF88DFFFE9800DFFFF81FFFFDFF4BFFFFF3),
    .INIT_08(256'hFC060103FFC00003FFFE0407FFE000103FFE00001FFFC0007FFC00000FFFE000),
    .INIT_09(256'h00203DFFC00023FC000203FFC00003FFF80003BFC000303FFC00021FFFD0007F),
    .INIT_0A(256'h027F8000200FE002007FFF80001BFC400200FF000003FFF400007FC000101FF8),
    .INIT_0B(256'h3C08000FFFE001043FA0000007C010007FFC800003F98002007E008007FFF800),
    .INIT_0C(256'h002081FF0008003880001FFF8002083FE0000003C20000FFEE001043FC000600),
    .INIT_0D(256'h8001000003FFE9A02200FE2008000800001FFFB000201FF8008003B00001FFF2),
    .INIT_0E(256'hCFFFFFC007F1C18033C00003FF3FFF0001FE0018005C00001FF8BFC1001FD300),
    .INIT_0F(256'h01A3027FC0007F9FA7FEFFEFD0700007F00003FEFEFFFCD87E040070BE00003F),
    .INIT_10(256'h0F9FFBBD07FFC700B807FFF800FC7FF3FC3C7DE005402FFC0007F1FB7F8D3FFF),
    .INIT_11(256'hFBF6FD01BFFFE01C7FFBDA03FD5F47C007FFFE00FBFFBFE07FBFFC4C007FFFC0),
    .INIT_12(256'hFFC23FFFFCC03FE5FFFE02FFFFFC3FFFFBF803FFCF7FC017FFFF01FFFFFF801F),
    .INIT_13(256'h25C03FFFE0FFFFFFED617F5C081F03FBBE03FFFFFF9FFFF44581FC3FFFE01FFF),
    .INIT_14(256'hFD400139FFE0F403005FDEE37FFFC207FFFF0E423003FFDEBFFFFFD9DFFFF1EC),
    .INIT_15(256'h00824013FF7F260000107E7FE03438047FDFFFD6800183FFFF05800087FFFF8F),
    .INIT_16(256'hE900001907FFFC0040000FFFBF800003B07FEFC0190C003FF7FA000003C7E3FE),
    .INIT_17(256'hFD90441000FFFBFC4000240FFFF80060041FFFFEC8000220FFF7C00008007FF3),
    .INIT_18(256'h7FF7C001B201FFFCC00A0002B7FFF83004300FFFE20041002BFFBFC0003880FF),
    .INIT_19(256'h1F183F830401FEFFDFC0230403FE83E011400BCFFCFC0818E01FFC0C0080023D),
    .INIT_1A(256'hA7FFFE7C03000000003FC208017FFFE3C0062003B001F001C013FFFFFC018000),
    .INIT_1B(256'h9FFCE803FF74003FBFFD1C4007FFCBC07FF28002FFFFE1C10054F2800BFC2141),
    .INIT_1C(256'h011BFBFFFA140207F00F2D1140003FFFFF800009FF4A68BFE80003FBFFD00000),
    .INIT_1D(256'hE8801C0003FFFFD01FFBFFFC0F0803E0000FFE3C31FFBFFF41E0203F00093CE0),
    .INIT_1E(256'hDFBFF3FFFFFF70BDBF100007FBFFFCFFFBFFF62FEE3CC0107E7DBF17FFBFFF01),
    .INIT_1F(256'hFFE1FDFE3E007FB3DF63FFFFFFFE3BFFE280DFFFFDFABFFFFFF607DBFED0007F),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n363,open_n364,addra[13]}),
    .dia({open_n368,open_n369,open_n370,open_n371,open_n372,open_n373,open_n374,1'b0,open_n375}),
    .rsta(rsta),
    .doa({open_n390,open_n391,open_n392,open_n393,open_n394,open_n395,open_n396,open_n397,inst_doa_i0_005}));
  // address_offset=0;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFF1FFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFF67EFE7FFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFC0FFFF80FFFFFFFFFFFFFFFFFF0FFFF87FFFFFFFFFFFFFFFFFF9FF),
    .INIT_02(256'h03FFFC007FFFFFFFFFFFFFFF807FFFC00FFFFFFFFFFFFFFFFC07FFFC03FFFFFF),
    .INIT_03(256'hFFFFFFFFFEFFC003FFFE007FFFFFFFFFFFFFFE003FFFE007FFFFFFFFFFD3FFF0),
    .INIT_04(256'hC0001FFFF81FFFFFFFFFFF7FFE0003FFFE00FFFFFFFFFFFFF7F8001FFFE00FEF),
    .INIT_05(256'hFFF1FFFFFFFFDCBF000FFFF83FFFEFFFFFFFFFF20000FFFF81FFF7FFFFFFEFFE),
    .INIT_06(256'hC079FFFFBFFFC7FE009FFFFF3F439FFFC7FFFC3FF81FFFFFFBFDDBFF00FFFFC3),
    .INIT_07(256'h0000018FFFFFC003F0FFFF0003FE000877FFFED81F0FFFF81FFE7C0087FFFFF3),
    .INIT_08(256'hFC05FE03FFC0000F800203FFFFE00FE03FFE00003800007EFFFC007F07FFE000),
    .INIT_09(256'h003FFE00407FF7FC0FFC01FFC000FFE00007FDFFC07FC03FFC0003FC00203F9F),
    .INIT_0A(256'hFC7FC7FFC00FE003FFFF80003FFFFC7FFC00FF000FFFF00C03FF7FC1FFC01FF8),
    .INIT_0B(256'h3C0FFFFFFE0003F83FBFFF8007C03FFFFFC3001FC3F87FFC007E00FFFFF81003),
    .INIT_0C(256'h000F81FCFFF00018FFFFFFFF4003F81FDFFF8003C3FFFFFFF0001FC3FFFFFC00),
    .INIT_0D(256'h0003FFFFFFFFCE201E01FC1FF0001FFFFFFFFF1000C01FC7FF0001BFFFFFFFF8),
    .INIT_0E(256'hCFE001800FE0BF000FFFFFFFFFBE000801FC0FE000BFFFFFFFFF8040C01FE0FF),
    .INIT_0F(256'h01C2FDFFFFFFFFFFA0029FEBE02E07FFFFFFFFFCFE0000DC7E03E03F7FFFFFFF),
    .INIT_10(256'hFFDFFB830007BE0007FBFFF7FFFCFFF00441FBE0043FDFFFFFFFF7FB800ABFBE),
    .INIT_11(256'h07F000FEFFFFEFFDFFFBC204027F803FFFFFFFFFF7FFBC00405DF803FFBFFFFF),
    .INIT_12(256'hFFFDFFFFFB000003FC01FDFFFFFFFBFFFBF800001F401FEFFFFFFFBFFFFE0020),
    .INIT_13(256'hD4003FC00F7FFFFFFD1FFFE3F02003FC00FFFFFFFFEFFFFDAB00043FC00FDFFF),
    .INIT_14(256'hFF3FFF83FFE003FE807FE00CFFFFFDF8FFFF11BDE003FC0047FFFFF6DFFFFA13),
    .INIT_15(256'h037DCFC3FF0037FFFFE381FFE00BC4F43FF001FE7FFE581FFF02FFFC07FE007F),
    .INIT_16(256'h0FFFFFE9F802FC00B787FFFF00FFFFFC3F801FC012B4FFFFF005FFFFFDF80FFE),
    .INIT_17(256'h01903BF03EFFFC1FBFFF83F00038005F07FFFFC0B7FFFC3F00078003F07FFFF8),
    .INIT_18(256'hFFC7FF7EB3FF00003FF3E03FFFFC7FDFFC3FF00015FFBF03DFFFC3BDFFD8FF00),
    .INIT_19(256'hE040007C0C01FFFFFFFFF907FC00001FE18017FFFCFFFFF0FFE00013FF3E01FF),
    .INIT_1A(256'h3FFFFF7FFDC1FFE000003C0000FFFFF3FFC63FFE00020FE0C00FFFFFFFFE807F),
    .INIT_1B(256'h7FF80004008FC03FFFFF0FC0FBFFC000000CFC03FFFFF3FF0FDBF0000001C080),
    .INIT_1C(256'hFE07FFFFF2D00FFFE00002C1BFE07FFFFF0600F6FF88004017FC07FFFFF0E00F),
    .INIT_1D(256'hE8FFFC00023FF83F1FFFFFF7EF0FFFE0001FFE43E1FFFFFF1DE0DFFE04026CE7),
    .INIT_1E(256'h1FC00FFFFFFEEFBDFFE8000003FC037FFFFFEFDFE1C38000007F80F7FFFFFFFF),
    .INIT_1F(256'h8FE9FFFF3F00007BE0C3FFFFFCFDBBFFF20080007E04FFFFFFCFB7DFFFC00040),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n423,open_n424,addra[13]}),
    .dia({open_n428,open_n429,open_n430,open_n431,open_n432,open_n433,open_n434,1'b0,open_n435}),
    .rsta(rsta),
    .doa({open_n450,open_n451,open_n452,open_n453,open_n454,open_n455,open_n456,open_n457,inst_doa_i0_006}));
  // address_offset=0;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h003FFFFFFFFFFFFFFFE00010000FFFFFFFFFFFFFFFFF98101FFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFC0003F000001FFFFFFFFFFFFFF0000F000007FFFFFFFFFFFFFF8000600),
    .INIT_02(256'hFC0000007FFFFFFFFFFE00007F8000000FFFFFFFFFFFF80003F8000003FFFFFF),
    .INIT_03(256'hFFFFFFFFFE003FFC0000007FFFFFFFFFFFC001FFC0000007FFFFFFFFFFD0000F),
    .INIT_04(256'h3FFFE000001FFFFFFFFFFF7FE1FFFC000100FFBFFFFFFFF7F007FFE000100FEF),
    .INIT_05(256'hFFF1FFFFFFFFDC00FFF000003FFFFFFFFFFFFFF1FFFF000001FFF7FFFFFFEFFE),
    .INIT_06(256'hC0000000400027FC009FFFFF3F4000003800003FF81BFFFFFBFFC000FF000003),
    .INIT_07(256'hFF00008FFFFFC000000000FFFC0E0008FBFFFED800000007E0007C000FFFFFF3),
    .INIT_08(256'hFC040000003FFFF0000007FFFFE000004001FFFFC00000FEFFFC000000001FFF),
    .INIT_09(256'hFFC00000007FF7FC000000003FFF00000007FEFFC000000003FFFC0000003FFF),
    .INIT_0A(256'hFE3FC00000001FFC000000003FEFFC40000000FFF000000403FF7FC000000007),
    .INIT_0B(256'h03F00000000003FC3F800000003FC0000000001FC3FC00000001FF0000001003),
    .INIT_0C(256'h000F81FF00000007000000004003F81FE00000003C00000000001FC1FC000400),
    .INIT_0D(256'h0001000000002FE00C00FFC0000000000000017001E00FF80000004000000000),
    .INIT_0E(256'h2FFFFF8007FF010003E00000007DFF0801FFF000001C00000003BFC0C01FFE00),
    .INIT_0F(256'hFE0200FFC000007FAFFD1FEFFFC00007F8000000FEFFF8FC7FFC00207F000000),
    .INIT_10(256'h001FFBBFF807BFFFC001FFF00002FFF7F380FBFFF8001FFE00000FFBFFF03FFF),
    .INIT_11(256'h03F700007FFFE0037FFBFDFC00DF7C2007FFFE0007FFBFFFC01FF7F0003FFFC0),
    .INIT_12(256'hFFE07FFFFF3FC003FC0001FFFFFC03FFFBF7FC003F80000FFFFF803FFFFFFFC0),
    .INIT_13(256'h1A003FC4007FFFFFFD3FFFBF03E003F80003FFFFFF8FFFFDE0FC043FC0103FFF),
    .INIT_14(256'hFF7FFC87FFEFF800007FE000FFFFFFE4FFFFFF004003FC000FFFFFFF5FFFFDF0),
    .INIT_15(256'hFF800037FF0037FFFFEF80FFFFB8080C3FE003FEFFFFB81FFFFF804007FE001F),
    .INIT_16(256'h06FFFFE7F800FFFF880007FF005FFFFFCF803FFFF804007FF007FFFFFE7807FF),
    .INIT_17(256'h03EF800000FFFC07FFFFBBF0003FFFC0000FFFC17FFFFDFF000FFFF500007FF8),
    .INIT_18(256'hFFC03F7F4DFF000480020001FFFC03FFFFCFF000080001001FFF803FFFF77F00),
    .INIT_19(256'hE0001F0000003FFFE03FFAFFFE0001E0010003FFFE03FFE73FE0021C0000001F),
    .INIT_1A(256'h3FFFFF43FDDFFFE0003F8000007FFFEC3FD9CFFE0003F8004007FFFF03FFFF7F),
    .INIT_1B(256'h80070007FF1FC01FFFFF03C0F80030007FE0F803FFFFF03F0F980E0003FE0180),
    .INIT_1C(256'hFE0FFFFFF2D00E001F800FF11FC03FFFFF0600F0007000FFFFFC03FFFFF0300F),
    .INIT_1D(256'hE88003FC023FE00E1FFFFFFFEF0C001FC00FFE83E0FFFFFFBFE0E001F800ECE8),
    .INIT_1E(256'h1C000FFFFFFFFFBD8007FE0003C0017FFFFFFFFFE0007FE0007C0077FFFFFFFE),
    .INIT_1F(256'hFFE9FE00C1F80000007FFFFFFFFFBBC00D7F800000017FFFFFFFFFDC003FF040),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n483,open_n484,addra[13]}),
    .dia({open_n488,open_n489,open_n490,open_n491,open_n492,open_n493,open_n494,1'b0,open_n495}),
    .rsta(rsta),
    .doa({open_n510,open_n511,open_n512,open_n513,open_n514,open_n515,open_n516,open_n517,inst_doa_i0_007}));
  // address_offset=0;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFF81FFFFFFFFFFFF83FFFFFFFFFC3FFFFFFFFFFFF8FFFFFFFFFFEFFFFF),
    .INIT_04(256'hFFFFFFFFFFE001FFFFFFFF801FFFFFFFFFFF007FFFFFFFF80FFFFFFFFFFFF01F),
    .INIT_05(256'h000FFFFFFFC0207FFFFFFFFFC0001FFFFFFC000FFFFFFFFFFE000FFFFFFFF001),
    .INIT_06(256'h400FFFFFFFFFF803FC9FFFFFC0407FFFFFFFFFC007DFFFFFFC01C7FFFFFFFFFC),
    .INIT_07(256'hFFFFFF8FFFFFE0000FFFFFFFFFF1FFF0FFFFFF1800FFFFFFFFFF83FF8FFFFFFC),
    .INIT_08(256'hFC0401FFFFFFFFFFFFFE07FFFFE0001FFFFFFFFFFFFFE0FEFFFC0000FFFFFFFF),
    .INIT_09(256'hFFFFFFFF807FF7FC0001FFFFFFFFFFFFFC07FEFFC0001FFFFFFFFFFFFFC03FFF),
    .INIT_0A(256'hFFFFC0003FFFFFFFFFFFFF003FE7FC4003FFFFFFFFFFFFFC03FFFFC0003FFFFF),
    .INIT_0B(256'hFFFFFFFFFFE003FFFF80007FFFFFFFFFFFFE001FFFFC0003FFFFFFFFFFFFE003),
    .INIT_0C(256'h000F7FFC0007FFFFFFFFFFFF8003F7FFC0007FFFFFFFFFFFFC001FBFF80003FF),
    .INIT_0D(256'hFFFCFFFFFFFFF7E00DFFFC000FFFFFFFFFFFFEF001FFFFC000FFFFFFFFFFFFF8),
    .INIT_0E(256'hF07FFFFFF7E000FFC01FFFFFFF87FF0FFEFE000FFF03FFFFFFFC3FC0FFEFC000),
    .INIT_0F(256'h001C00003FFFFFC02FFE0FEFE001F80007FFFFFD06FFF0C3FE001FC000FFFFFF),
    .INIT_10(256'hFFE003FE0007BF000000000FFFFF0077F800FFF003000001FFFFF0037FC03FFE),
    .INIT_11(256'h01F8FE0000001FFF8003F800005F03C0000001FFF8003FC0401DF00C0000003F),
    .INIT_12(256'h001F000079400003FBFE00000003FC0003E000003FBFE00000007FC0007F0000),
    .INIT_13(256'h00003FC3F000000002FFFFC0042003FCFF000000007000041100043FDFF00000),
    .INIT_14(256'h00FFFF07FFEF0000007FE0F000001FE8FFFFE0000003FC1F000000079FFFFE00),
    .INIT_15(256'hFC000013FF008FFFFFEC00FFFFC000043FE01800FFFFE01FFFF8804007FE0380),
    .INIT_16(256'h07FFFFEE0000FFFF080007FF007FFFFFF0003FFFE004003FF003FFFFFF8007FF),
    .INIT_17(256'h01FFFC0000FFFC07FFFFFC00003FFFC0000FFFC07FFFFDC00007FFF800007FF8),
    .INIT_18(256'hFFC03F7FFE0000037FFC0001FFFC03FFFFF000000FFFC1001FFFC03FFFFF8000),
    .INIT_19(256'h007FE0FFF0003FFFE03FFBF80000FE1FFF0003FFFE03FFFFC00001E3FFE0001F),
    .INIT_1A(256'h3FFFFF83FA3E001FFFC07FF8007FFFF03FDFF0003FFC07FF4007FFFE03FFFF80),
    .INIT_1B(256'h0007FFF800E0003FFFFFF3FF00003FFF801F0002FFFFFE3FF06003FFFC03FE00),
    .INIT_1C(256'h0007FFFFFDEFF0000FFFF00E80007FFFFFF9FF0000FFFF00000003FFFFFFBFF0),
    .INIT_1D(256'h170003FFFDC018001FFFFFFFF0F0001FFFF0018000FFFFFFFE1F0001FFFF3318),
    .INIT_1E(256'hE3C007FFFFFFFF420007FFFFFC3C007FFFFFFFF018003FFFFF838007FFFFFFFF),
    .INIT_1F(256'hFFEE000001FFFFFBC07FFFFFFFFFC400007F7FFFFC01FFFFFFFFF820001FFFBF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_008 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n543,open_n544,addra[13]}),
    .dia({open_n548,open_n549,open_n550,open_n551,open_n552,open_n553,open_n554,1'b0,open_n555}),
    .rsta(rsta),
    .doa({open_n570,open_n571,open_n572,open_n573,open_n574,open_n575,open_n576,open_n577,inst_doa_i0_008}));
  // address_offset=0;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hBFFFFFFFFFFFFFFFFC7FFFFFFFBFFFFFFFFFFFFFFFD3FFFFFFFE3FFFFFFFFFFF),
    .INIT_07(256'hFFFFFF803FFFFFFFFFFFFFFFFFFFFFF807FFFFE7FFFFFFFFFFFFFFFF80FFFFFF),
    .INIT_08(256'hFFFBFFFFFFFFFFFFFFFE0007FFDFFFFFFFFFFFFFFFFFF081FFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFF80400FFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFC0403F),
    .INIT_0A(256'h01FFFFFFFFFFFFFFFFFFFF00001FFFBFFFFFFFFFFFFFFFFC0000FFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFE00203FFFFFFFFFFFFFFFFFFFE00203FFFFFFFFFFFFFFFFFFFF000),
    .INIT_0C(256'h0010FFFCFFFFFFFFFFFFFFFFC0020FFFDFFFFFFFFFFFFFFFFC00007DFBFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFE3E003FFFC3FFFFFFFFFFFFFFF70011FFFC7FFFFFFFFFFFFFFF8),
    .INIT_0E(256'hF01FFF7FFFE07FFFFFFFFFFFFF81FF07FFFE0FFFFFFFFFFFFFFC7FC03FFFC1FF),
    .INIT_0F(256'h00FFFFFFFFFFFF805FFF9017E01FFFFFFFFFFFFE01FFFB3FFE03FFFFFFFFFFFF),
    .INIT_10(256'hFFC0047FF8007F003FFFFFFFFFFE000FFF8107F007FFFFFFFFFFF004FFF8407E),
    .INIT_11(256'h03F001FFFFFFFFFF00043FFC00BF001FFFFFFFFFF80043FFC003F003FFFFFFFF),
    .INIT_12(256'hFFFF8000017FC003F801FFFFFFFFFC00041FFC003F801FFFFFFFFFE00001FFC0),
    .INIT_13(256'h1E003FC00FFFFFFFFC00000007E003FC00FFFFFFFFE0000201FC043FC00FFFFF),
    .INIT_14(256'hFF80000000100000007FE00FFFFFE000000000006003FC00FFFFFFF800000000),
    .INIT_15(256'h0001FFF3FF0078000000000000000FFC3FE007FF000000000000807C07FE007F),
    .INIT_16(256'h06000000000100000FFFFFFF0040000000000000003BFFFFF000000000000000),
    .INIT_17(256'h000003FFFFFFFC07800000000000007FFFFFFFC07000020000000001FFFFFFF8),
    .INIT_18(256'hFFC03F80000000000001FFFFFFFC03E00000000000003EFFFFFFC03C00100000),
    .INIT_19(256'h000000000FFFFFFFE03FC4000000000000FFFFFFFE03F81000000000001FFFFF),
    .INIT_1A(256'hCFFFFE03FC00000000000007FFFFFFE03FC0000000000000BFFFFFFF03FE0000),
    .INIT_1B(256'h00000000001FFFDFFFFF03C00000000000007FFDFFFFF03F00000000000001FF),
    .INIT_1C(256'hFFFFFFFFF0C000000000000FFFFFFFFFFF0000000000000007FFFFFFFFF03000),
    .INIT_1D(256'h0000000001FFE7FFFFFFFFFFE0000000001FFF7FFFFFFFFF3E00000000001FF7),
    .INIT_1E(256'hFC3FFFFFFFFFFF0000000003FFC3FFFFFFFFFFF0000000003FFE7FFBFFFFFFFF),
    .INIT_1F(256'hFFE800000000FFC43F8FFFFFFFFF8000000007FF83FEFFFFFFFFF8000000007F),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n603,open_n604,addra[13]}),
    .dia({open_n608,open_n609,open_n610,open_n611,open_n612,open_n613,open_n614,1'b0,open_n615}),
    .rsta(rsta),
    .doa({open_n630,open_n631,open_n632,open_n633,open_n634,open_n635,open_n636,open_n637,inst_doa_i0_009}));
  // address_offset=0;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFF701FFFFFFFFFFFFFFFFFFFFFFF07FFFFFFFFFFFFFFFFFFFFFFF0FFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFF8007FFFFFFFFFFFFFFFFFFFFF800FFFFFFFFFFFFFFFFFFFFFF803F),
    .INIT_0A(256'h003FFFFFFFFFFFFFFFFFFFFFC007FFFFFFFFFFFFFFFFFFFBFC007FFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFC),
    .INIT_0C(256'hFFE001FFFFFFFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFE003FFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFE01FF000FFFFFFFFFFFFFFFFFF0FFE001FFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hF00000000FFFFFFFFFFFFFFFFF8000F000FFFFFFFFFFFFFFFFFC003F000FFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFF8000006007FFFFFFFFFFFFFFFE000004007FFFFFFFFFFFFFFF),
    .INIT_10(256'hFFC0000007F83FFFFFFFFFFFFFFE0000007E07FFFFFFFFFFFFFFF0000007807F),
    .INIT_11(256'hFFFFFFFFFFFFFFFF00000003FF3FFFFFFFFFFFFFF80000003FE3FFFFFFFFFFFF),
    .INIT_12(256'hFFFF800000803FFFFFFFFFFFFFFFFC00000003FFFFFFFFFFFFFFFFE00000003F),
    .INIT_13(256'hE1FFFFFFFFFFFFFFFC000000F81FFFFFFFFFFFFFFFE000000E03FBFFBFFFFFFF),
    .INIT_14(256'hFFFFFC0000000FFFFFBFFFFFFFFFFFF0000000FF9FFFFFFFFFFFFFFF8000000F),
    .INIT_15(256'h007E000FFFFFFFFFFFF000000007F003FFFFFFFFFFFF800000007F83FBFFFFFF),
    .INIT_16(256'hF9FFFFF000000000700007FFFFBFFFFF8000000007C0007FFFFFFFFFFC000000),
    .INIT_17(256'h0000000000FFFBF87FFF800000000000000FFFBF8FFFFC000000000600007FFF),
    .INIT_18(256'hFFFFC0FF8000000000000001FFFFFC1FFC000000000000001FFFFFC3FFE00000),
    .INIT_19(256'h0000000000003FFFFFC03C0000000000000003FFFFFC07E0000000000000003F),
    .INIT_1A(256'h0FFFFE3C0000000000000000007FFFE7C0200000000000000007FFFEFC018000),
    .INIT_1B(256'h000000000000001FFFFF0C000000000000000000FFFFF1C00000000000000000),
    .INIT_1C(256'h000FFFFFF00000000000000000007FFFFF00000000000000000003FFFFF04000),
    .INIT_1D(256'h00000000000000001FFFFFF8000000000000000000FFFFFF0000000000000000),
    .INIT_1E(256'h00000FFFFFFFF000000000000000007FFFFFFE000000000000000003FFFFFFC0),
    .INIT_1F(256'hFFF00000000000000003FFFFFFFC00000000000000007FFFFFFF800000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n663,open_n664,addra[13]}),
    .dia({open_n668,open_n669,open_n670,open_n671,open_n672,open_n673,open_n674,1'b0,open_n675}),
    .rsta(rsta),
    .doa({open_n690,open_n691,open_n692,open_n693,open_n694,open_n695,open_n696,open_n697,inst_doa_i0_010}));
  // address_offset=0;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFE7FFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFF83FFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFC003FFFFFFFFFFFFFFFFFFFFFC00FFFFFFFFFFFFFFFFFFFFFF803FFFFFF),
    .INIT_03(256'hFFFFFFFF80FFFFFFFFFE000FFFFFFFFFFC3FFFFFFFFFE006FFFFFFFFFFF7FFFF),
    .INIT_04(256'hDFFFFFFFF80003FFFFFFFF001FFFFFFFFF01007FFFFFFFF807FFFFFFFFE0000F),
    .INIT_05(256'h0015FFFFFFC0CEBFFFFFFFF800001FFFFFFC0193FFFFFFFF800007FFFFFFF002),
    .INIT_06(256'hF3F5FFFFFFFFC403FA8FFFFF3B7F9FFFFFFFFC0007EFFFFFF80AD9FFFFFFFFC0),
    .INIT_07(256'hFFFFFFB85FFFFFFFF1FFFFFFFFF3FFFB07FFFE5FFF4FFFFFFFFE41FF3BFFFFF3),
    .INIT_08(256'hFFFFFE03FFFFFFFFBFFFFC06FFFFEFF03FFFFFFFFFFFFF807FFCFF3E17FFFFFF),
    .INIT_09(256'hFFFFFFFFFFC02FFFFFFC01FFFFFFFFFFFBFA03FFFFFFE03FFFFFFFFFFFFF807F),
    .INIT_0A(256'h023FF7FFC00FFFFFFFFFFF7F8017FFBFFC02FF7FFFFFFFF3F801FFFFFFE01FFF),
    .INIT_0B(256'h3FFFFFFFFDFFFF041FFFFFC007FFFFFFFFFCFFC003FFFFFC007FFFFFFFFFFFFE),
    .INIT_0C(256'hFFF101FCFFF0001FFFFFFFFF9FFD181FFFFFC003FFFFFFFFFDFFD083FFFFFC00),
    .INIT_0D(256'h000FFFFFFFFFFC3FF201FDBFF8001FFFFFFFFF17FD201FC7FF0001FFFFFFFFF7),
    .INIT_0E(256'hCF9001B80FFEFE007FDFFFFFFFB800F801FFCFF000FFFFFFFFFAA07F0007DFFF),
    .INIT_0F(256'hFE41FFFFFFFFFFDFD0026403EFBE07FBFBFFFFFEF9002604FCFBE00FFFFFFFFF),
    .INIT_10(256'hFFFFF80107F83EFF9FFDFFF7FFFFFFD4007F07EFF47FDFFFFFFFF9FD0107C07F),
    .INIT_11(256'hFBFDFFFF7FFFFFFDFFF82603FF4FF9DFFFFFFFFFFFFF8400FFE1F3A5FFBFFFFF),
    .INIT_12(256'hFFFDBFFF91003FFBFFFEFFFFFFFDFFFFF82803FFBF3FFFE7FFFFFFFFFFC0803F),
    .INIT_13(256'hC1FFFFFFFFBFFFFFFB1FBFC0F83FFFFFFFFBFFFFFFFFFFFC0A83FBFFFFFFDFFF),
    .INIT_14(256'hFD400539FFE18BFDFFFFFFEF7FFFE21B7FFF003F9FFFFFFEFBFFFDDD3FFFF803),
    .INIT_15(256'h007F8013FF7FB40000127F7FE00FC503FFEFDFFE800007FFFF043FC67BFFFF7F),
    .INIT_16(256'hE50000101FFCFC007D080BFFBFE00003107FCFC022AC007FF7FE00000417E7FE),
    .INIT_17(256'hFC9187C040FFFBE38000A00FFFB800378417FFBE700004007FFF800374007FFB),
    .INIT_18(256'hFFF03F804001FFF9C009C001FFFFC7E012000FFFE4001F001FFFBC7E003001FF),
    .INIT_19(256'h3FBFE1030001BFFFD03FE60401FE7F3011C00DFFFE03F028200FFEF4007C003F),
    .INIT_1A(256'h5FFFFF43F942000FFFE0030000BFFFC43FE800038FFE0800C007FFFE03FE8000),
    .INIT_1B(256'h0000FFF803003FFFFFFF12C000008C7F803047FEFFFFF33E01870D7FFA00017E),
    .INIT_1C(256'h02EFFFFFFCD80004107E4C96C03F3FFFFF8A000000CFDF80C803FBFFFFE0A800),
    .INIT_1D(256'hF4000401FE3FF401DFFFFFFBFE0000003FFFFE000EFFFFFFDFE0000207FD4BE8),
    .INIT_1E(256'h1FC00FFFFFFEFF7E7FF000F807FC007FFFFFEFDFF000001FE07D8009FFFFFFFD),
    .INIT_1F(256'h8FEFC3FFFE838037C075FFFFFCFDFE3FFEC070003C01FFFFFFCFBFF7FFC01F80),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_011 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n723,open_n724,addra[13]}),
    .dia({open_n728,open_n729,open_n730,open_n731,open_n732,open_n733,open_n734,1'b0,open_n735}),
    .rsta(rsta),
    .doa({open_n750,open_n751,open_n752,open_n753,open_n754,open_n755,open_n756,open_n757,inst_doa_i0_011}));
  // address_offset=0;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h003FFFFFFFFFFFFFFFE00000000FFFFFFFFFFFFFFFFF18001FFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFC00000000001FFFFFFFFFFFFFF00000000007FFFFFFFFFFFFFF8000000),
    .INIT_02(256'h000000003FFFFFFFFFFE0000000000000FFFFFFFFFFFF8000000000003FFFFFF),
    .INIT_03(256'hFFFFFFFF800000000000000FFFFFFFFFFC00000000000006FFFFFFFFFFC00000),
    .INIT_04(256'h20000000000003FFFFFFFF00000000000000003FFFFFFFF0000000000010000F),
    .INIT_05(256'h0012FFFFFFC003800000000000001FFFFFFC000800000000000007FFFFFFE000),
    .INIT_06(256'h3FF8000000002400051FFFFF00FF8000000000000017FFFFF801F80000000000),
    .INIT_07(256'h0000004FBFFFDFFFF00000000002000C7FFFFE3FFF0000000000400044FFFFF0),
    .INIT_08(256'hFFFFFE0000000000000203FFFFFFFFE0400000000000007CFFFFFFFF00000000),
    .INIT_09(256'h00000000007FDFFFFFFE0000000000000401FDFFFFFFE0000000000000007FFF),
    .INIT_0A(256'hFDFFFFFFC0000000000000807FFFFFFFFC0000800000000C07FE7FFFFFC00000),
    .INIT_0B(256'h00000000022000FBFFBFFF80000000000000001FFFFFFFFC0000000000000001),
    .INIT_0C(256'h000EFDFCFFF80000000000006000E7DFDFFF80000000000000000F7FFBFFF800),
    .INIT_0D(256'h0001000000001C001FFEFC3FF00000000000018802DFFFC7FF0000000000000C),
    .INIT_0E(256'h3F8000C7FFE0FE0003E0000000FA0007FFFE0FF0001C000000048000FFFFC1FF),
    .INIT_0F(256'h006000FFC000001F8001EFFFE03E0007F8000003F80015DB7E03E0107F000000),
    .INIT_10(256'h003FF840FFFFBF002003FFF00003FFC00FFFFDF006003FFE000005F8807FBFFF),
    .INIT_11(256'hFFF00000FFFFF0017FF803FFFFFF820007FFFE0007FF801F7FFFF00A007FFFC0),
    .INIT_12(256'hFFE2FFFF86BFFFFFF80101FFFFFC07FFF807FFFFFF80001FFFFF805FFFC27FFF),
    .INIT_13(256'h2DFFFFC4007FFFFFF93FBFBF03FFFFF80007FFFFFFAFFFFDF5FFFFFF80103FFF),
    .INIT_14(256'hFF400639FFEE7C03FFFFE010FFFFE20BFFFFFFC03FFFFC010FFFFFFCBFFFFDFC),
    .INIT_15(256'hFF803FFBFF80340000007EFFFFB033FFBFF023FE800007DFFFFBC03BFFFE009F),
    .INIT_16(256'h130000000FFDFFFF807FF7FF40A00000907FEFFFD947FFFFF80200000607E7FF),
    .INIT_17(256'hFCEE000FFEFFF8040000200FFFBFFF80FBEFFF80000004007FFFFFF50FFF7FFC),
    .INIT_18(256'hFFC800004000FFFCC0061FFFFFFC440012000FFFE00041FFFFFFC042002000FF),
    .INIT_19(256'h1F801F00F3FE7FFFF000060401FE01E00F3FFBFFFF000838200FFC1C00E3FDFF),
    .INIT_1A(256'h7FFFFF0000200000003FC1FFFFFFFFFC000800018003F01F7FEFFFFF00008000),
    .INIT_1B(256'h7FFF0807FF7FC01FFFFF114007FF60007FF3F800FFFFF300000FF20003FC3F80),
    .INIT_1C(256'hFC0FFFFFF48001FBFF800FF9DFC07FFFFF8E000FFFB800FFFFFC03FFFFF09800),
    .INIT_1D(256'h087FFBFE01C01C0E3FFFFFFC0103FFFFC0000183E1FFFFFF60001FFDFC00D418),
    .INIT_1E(256'hE3C00FFFFFFFF001FFFFFF07F83C017FFFFFFF200FFFBFE01F83C073FFFFFFC2),
    .INIT_1F(256'hFFF43DFFFFF87FFFC077FFFFFFFE01FFFEBF8FFFBC017FFFFFFF800BFFDFE03F),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_012 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n783,open_n784,addra[13]}),
    .dia({open_n788,open_n789,open_n790,open_n791,open_n792,open_n793,open_n794,1'b0,open_n795}),
    .rsta(rsta),
    .doa({open_n810,open_n811,open_n812,open_n813,open_n814,open_n815,open_n816,open_n817,inst_doa_i0_012}));
  // address_offset=0;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFEEFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'h800FFFFFFFFFFBFFFF1FFFFFFF007FFFFFFFFFFFFFF3FFFFFFFE07FFFFFFFFFF),
    .INIT_07(256'hFFFFFFF81FFFE0000FFFFFFFFFFDFFFF07FFFFC000FFFFFFFFFFBFFFF0FFFFFF),
    .INIT_08(256'hFC0001FFFFFFFFFFFFFDF807FFC0001FFFFFFFFFFFFFFF80FFFC0000FFFFFFFF),
    .INIT_09(256'hFFFFFFFFBFC00FFC0001FFFFFFFFFFFFFFF800FFC0001FFFFFFFFFFFFFDF803F),
    .INIT_0A(256'h01BFC0003FFFFFFFFFFFFF7FC00FFC0003FFFFFFFFFFFFFFFC00FFC0003FFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFE03FF80007FFFFFFFFFFFFFFFC03FFC0003FFFFFFFFFFFFFFFC),
    .INIT_0C(256'hFFE0FFFF0007FFFFFFFFFFFFFFFE0FFFE0007FFFFFFFFFFFFFFFE07FFC0007FF),
    .INIT_0D(256'hFFFCFFFFFFFFE7FFF1FEFFC00FFFFFFFFFFFFE7FFF1FFFF800FFFFFFFFFFFFFF),
    .INIT_0E(256'hF01FFFFFFFFF01FFC01FFFFFFF83FFF7FFFFF00FFF03FFFFFFFF3FFF3FFFFE00),
    .INIT_0F(256'hFF9E00003FFFFFE00FFFF007FFC1F80007FFFFFE00FFFC3FFFFC1FE000FFFFFF),
    .INIT_10(256'hFFC0003FFFF83FFFC000000FFFFD0047FFFE07FFFB000001FFFFFA007FFF807E),
    .INIT_11(256'hFFFFFE0000000FFF80003FFFFF1F7FE0000001FFF80003FFFFE1FFFC0000003F),
    .INIT_12(256'h001F800001FFFFFFFFFE00000003FC00001FFFFFFFFFE00000007FE00041FFFF),
    .INIT_13(256'hFFFFFFC3F000000004FFBFC0FFFFFFFCFF000000004000040FFFFFFF9FF00000),
    .INIT_14(256'h00C00645FFEF0FFFFFFFE0F000000218FFFFE0FFFFFFFC1F000000049FFFFE0F),
    .INIT_15(256'hFC7FF01FFF008C00001001FFFFC7FF07FFE018008000003FFFF8FFC3FFFE0380),
    .INIT_16(256'h090000100803FFFF7FF807FF0020000010002FFFE7FF007FF006000006001FFF),
    .INIT_17(256'h02FFFFFFC0FFF81800002000007FFFFFF80FFF8180000400800FFFFEF780FFF8),
    .INIT_18(256'hFFC7C00040000004BFFFFFC1FFFC3800120000001FFFFFFC1FFFC38200300000),
    .INIT_19(256'h00001FFFFFFE7FFFEFC00604000101FFFEFFE3FFFEFC00282010021FFFFDFC3F),
    .INIT_1A(256'h7FFFFF7C03E00000003FBFFFFF7FFFF3C01800004003F7FFFFE7FFFEFC000000),
    .INIT_1B(256'h8000F807FFE0003FFFFF1C3FF8000C007FEF8000FFFFF2C1FF88010003FFFE00),
    .INIT_1C(256'h000FFFFFFCFFFE00007F0FF040007FFFFF8DFFF0008FC0FFF80003FFFFF0C7FF),
    .INIT_1D(256'hFF800003FE0004001FFFFFFFFFFC00003FE0000001FFFFFFFFFFE00007FCE000),
    .INIT_1E(256'h00000FFFFFFFFFFF800001FC0000007FFFFFFFFFF800401FC0004003FFFFFFFF),
    .INIT_1F(256'hFFFBFE0000070004007BFFFFFFFFFFC00100F8004001FFFFFFFFFFFC00200F80),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_013 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n843,open_n844,addra[13]}),
    .dia({open_n848,open_n849,open_n850,open_n851,open_n852,open_n853,open_n854,1'b0,open_n855}),
    .rsta(rsta),
    .doa({open_n870,open_n871,open_n872,open_n873,open_n874,open_n875,open_n876,open_n877,inst_doa_i0_013}));
  // address_offset=0;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFE3FFFFFFFC3FFFFFFFFFFFFFFF7FFFFFFFC7FFFFFFFFFFFFFFFF),
    .INIT_0E(256'hF07FFF7FFFE07FFFFFFFFFFFFF85FFFFFFFE0FFFFFFFFFFFFFFC7FFFFFFFC1FF),
    .INIT_0F(256'h00FFFFFFFFFFFFC07FFFFFFFE01FFFFFFFFFFFFE07FFFFFFFE03FFFFFFFFFFFF),
    .INIT_10(256'hFFC007FFFFFFFF003FFFFFFFFFFF003FFFFFFFF007FFFFFFFFFFF807FFFFFFFE),
    .INIT_11(256'hFFF001FFFFFFFFFF0007FFFFFFFF001FFFFFFFFFF8007FFFFFFFF003FFFFFFFF),
    .INIT_12(256'hFFFF800079FFFFFFF801FFFFFFFFFC0007FFFFFFFF801FFFFFFFFFE0003FFFFF),
    .INIT_13(256'hFFFFFFC00FFFFFFFFC004000FFFFFFFC00FFFFFFFFE000020FFFFFFF800FFFFF),
    .INIT_14(256'hFFBFFA7A00100FFFFFFFE00FFFFFFDEB000000FFFFFFFC00FFFFFFFB2000000F),
    .INIT_15(256'h007FCFFFFF007BFFFFE07F000007FCFFFFE007FF7FFF87E00000FFFFFFFE007F),
    .INIT_16(256'h00FFFFE00FFE00007F87FFFF001FFFFF907FD00007F8FFFFF001FFFFFA07F800),
    .INIT_17(256'hFF0003F03FFFF8007FFFA00FFFC0007F07FFFF800FFFF800FFF80007F87F7FF8),
    .INIT_18(256'hFFC000FFC000FFFC8001E03FFFFC001FEE000FFFF0003E03FFFFC001FFC000FF),
    .INIT_19(256'h1F801F000C01BFFFE0003A0401FF01E001C01FFFFE0007C8201FFE1C001E03FF),
    .INIT_1A(256'h8FFFFF4003E00000003F800000FFFFF800180001C003F000801FFFFE00018000),
    .INIT_1B(256'hFFF8F807FF1FFFDFFFFF103FFFFFCC007FE07FFFFFFFF200FF8FFD0003FC01FF),
    .INIT_1C(256'hFFFFFFFFFC3FFFFFF07F0FFFBFFFFFFFFF8FFFFFFF8FC0FFFFFFFFFFFFF08FFF),
    .INIT_1D(256'hFFFFFC03FFFFE3FFFFFFFFF81FFFFFE03FFFFF7FFEFFFFFFC1FFFFFE07FCDFF7),
    .INIT_1E(256'hFC3FFFFFFFFFF0FFFFF801FFFFC3FFFFFFFFFE0FFFFFC01FFFFE3FFFFFFFFFC0),
    .INIT_1F(256'hFFE7FFFFFE07FFC03F8FFFFFFFFC7FFFFF80FFFF83FEFFFFFFFF87FFFFE00FFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_014 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n903,open_n904,addra[13]}),
    .dia({open_n908,open_n909,open_n910,open_n911,open_n912,open_n913,open_n914,1'b0,open_n915}),
    .rsta(rsta),
    .doa({open_n930,open_n931,open_n932,open_n933,open_n934,open_n935,open_n936,open_n937,inst_doa_i0_014}));
  // address_offset=0;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFD87FFFFFFFFFFFFFFFFFFFFFFF4FFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFF80FFFFFFFFFFFFFFFFFFFFFFF81FFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFF001FFFFFFFFFFFFFFFFFFFFEF803FFFFFFFFFFFFFFFFFFFFDF807FF),
    .INIT_17(256'h01FFFFFFFFFFFFFFFFFFDFF0003FFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFBFFF00037FFFFFFFFFFFFFFFFDFFF0000FFFFFFFFFFFFFFFFFFFFF00),
    .INIT_19(256'hE07FE0FFFFFFFFFFFFFFFDFBFE00FE1FFFFFFFFFFFFFFFF7DFE001E3FFFFFFFF),
    .INIT_1A(256'hFFFFFEBFFC1FFFFFFFC07FFFFFFFFFE7FFE7FFFE3FFC0FFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h000707F800FFFFFFFFFFEFC0000033FF801FFFFFFFFFFDFF007002FFFC03FFFF),
    .INIT_1C(256'hFFFFFFFFF3C000000F80F00FFFFFFFFFFF70000000703F0007FFFFFFFFFF7000),
    .INIT_1D(256'h000003FC01FFFFFFFFFFFFFFE000001FC01FFFFFFFFFFFFF3E000001F8033FFF),
    .INIT_1E(256'hFFFFFFFFFFFFFF000007FE03FFFFFFFFFFFFFFF000003FE03FFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFF8000001F8FFFFFFFFFFFFFFFF8000007F07FFFFFFFFFFFFFFF800001FF07F),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_000000_015 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n963,open_n964,addra[13]}),
    .dia({open_n968,open_n969,open_n970,open_n971,open_n972,open_n973,open_n974,1'b0,open_n975}),
    .rsta(rsta),
    .doa({open_n990,open_n991,open_n992,open_n993,open_n994,open_n995,open_n996,open_n997,inst_doa_i0_015}));
  // address_offset=8192;data_offset=0;depth=1508;width=4;num_section=1;width_per_section=4;section_size=16;working_depth=2048;working_width=4;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("4"),
    .DATA_WIDTH_B("4"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h111105555221899999533333555333666665333288CFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h2223887DFFFFFFFFFFFFFFFFFFFFFEEEFFFFFFFFFE2332222220111111111111),
    .INIT_02(256'hFFFFF0222222222211111111111111111111552989A233333332555633666752),
    .INIT_03(256'h101442333333333655555366732222288898FFFFFFFFFFFFFFFFFFFFEEEEFFFF),
    .INIT_04(256'hBEFFFFFFFFFFFFFFFFFEEEEEFFFFFFFFFFF22222222201111111111111111112),
    .INIT_05(256'h1222222230111111111333333333336333333333332555555365322222288887),
    .INIT_06(256'h3333335555555652222222288889ACFFFFFFFFFFFFFFFFFEEEEEFFFFFFFFFFDC),
    .INIT_07(256'hFFFFFFFFFFEEEEEEFFFFFFFFCCCCCA1121222011101111443333333333663333),
    .INIT_08(256'h2211111123444233333335666333333332555555376B22222228888AAAEFFFFF),
    .INIT_09(256'h5467777752222228985AAAACFFFFFFFFFFFFFFEEEEEEFFFFFFDCCCCCCCCA1122),
    .INIT_0A(256'hFEEEEEEEFFFFECCCCCCCCCCCCA22220111133444433333333666664333333555),
    .INIT_0B(256'h4444443333333666666333332564767677777623228998AAAAAACFFFFFFFFFFF),
    .INIT_0C(256'h777422998AAAAAAA9CFFFFFEFFFFEEEEEEEEFFFCCCCCCCCCCCCCCCCA31311143),
    .INIT_0D(256'hFCCCCCCCCCCCCCCCCCCDCC200344444444443333566666663233554676777777),
    .INIT_0E(256'h33336666666663334C6777777777777772B9AAAAAAAAAACFFFFEFFFFEEEEEEEE),
    .INIT_0F(256'hAAAAAAAAAAADFFFEFFFEEEEEEEECCCCCCCCCCCCCCCCCCCCCCCB7643443444444),
    .INIT_10(256'hCCCCCCCCB8899998989A844444444333666666666737766777777777777765AA),
    .INIT_11(256'h667A00233479999999999999999999AAAAAAAAAACFFFFFFEEEEEECCCCCCCCCCC),
    .INIT_12(256'hAAAAACFFFFEEEEECCCCCCCCCCCBCCD9999999999999999999999974333276666),
    .INIT_13(256'h99999899999888898898977FD0002344444555566677788899999999999999AA),
    .INIT_14(256'h88888999999A9AAABABBBA9999AAAAAAAAEFFFEEECCCCCCCCBBC989999999999),
    .INIT_15(256'hFEECCCCCCA899999999999999999999998887766666655544566555566666777),
    .INIT_16(256'h999889987777778777888888999999999AAAAABBBBBBBCBBCCCDDDDDDEDBAAAC),
    .INIT_17(256'h0000000000000000000000000000ECCA889899CCCDCCCCCCBBBBBBBBA9AAA999),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_008192_000 (
    .addra({addra[10:0],2'b11}),
    .clka(clka),
    .csa(addra[13:11]),
    .dia({open_n1026,open_n1027,open_n1028,open_n1029,open_n1030,4'b0000}),
    .rsta(rsta),
    .doa({open_n1045,open_n1046,open_n1047,open_n1048,open_n1049,inst_doa_i4_003,inst_doa_i4_002,inst_doa_i4_001,inst_doa_i4_000}));
  // address_offset=8192;data_offset=4;depth=1508;width=4;num_section=1;width_per_section=4;section_size=16;working_depth=2048;working_width=4;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("4"),
    .DATA_WIDTH_B("4"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h666664888E0E222222246666202666422222888A880FFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h8880886DFFFFFFFFFFFFFFFFFFFFDBBBDFFFFFFF0C0EEEEEEEE4666666668866),
    .INIT_02(256'hFFFFF70EEEEEEEEC6666666888666666664A88022244666666660000662244E8),
    .INIT_03(256'h64E0A488666666600000C6224A8888848868FFFFFFFFFFFFFFFFFFFFBBBBDFFF),
    .INIT_04(256'hA9FFFFFFFFFFFFFFFFFBBBBBFFFFFFFFFF4EEEEEEEEE46666668886666666666),
    .INIT_05(256'hAEEEEEEEE466668888800000000000E486666666662000000642A88888868888),
    .INIT_06(256'h666668200000020888888868888685FFFFFFFFFFFFFFFFFBBBBBFFFFFFFFFD57),
    .INIT_07(256'hFFFFFFFFFFBBBBBBFFFFFFFF35555FECECEEE466668886220000000000EE8666),
    .INIT_08(256'hEA66668882222000000006CCC68666666400000031F6888888A88888BBBFFFFF),
    .INIT_09(256'h22C31FF1BA8888A888BBBBB5FFFFFFFFFFFFFDBBBBBBFFFFFF535555535DAEEE),
    .INIT_0A(256'hFBBBBBBBFFFFB5555555555533CCEE6668822222220000000EEEEE6666666000),
    .INIT_0B(256'h2222222000000CEEEEC8666642E24DF11F11FFE88886A7BBBBBB5FFFFFFFFFFF),
    .INIT_0C(256'hFF1A8888B9BBBBBBB5FFFFFDFFFFBBBBBBBBFDF5555555555555555F0EE66822),
    .INIT_0D(256'hF335555555555555555337C442222222222200008EEEEECC686800CFFFFFFFFF),
    .INIT_0E(256'h2000CEEEEEEEC686061FFFFFFFFFFFFF4C09BBBBBBBBBB5FFFFDFFFFBBBBBBBB),
    .INIT_0F(256'hBBBBBBBBBBB5FFFDFFFBBBBBBBD3333333333333333333333311C40022222222),
    .INIT_10(256'h33333333F35777797779342222222000EEEEEEEECC661F1FFFFFFFFFFFFF1FBB),
    .INIT_11(256'hCE0279F3353BBBBBDBBBBBBBBBBBBBBBBBBBBBBB3FFDFFFBBBBBB13333333333),
    .INIT_12(256'hBBBBB5FFFFBBBBB333333333331337777777777777777777777955424EEECECC),
    .INIT_13(256'h777777777777775977777574C7FB15135579BBDFFF1335579BBBBBBBBBBBBBBB),
    .INIT_14(256'h5579799999BDBDBDFF111FBBBBBBBBBBBB9FFDBBD33333333113757777777777),
    .INIT_15(256'hFBB333333D57777777777777777777797775131DBDBD9BB997DD9DFDDFFF1135),
    .INIT_16(256'h99975533355533113555379979999BBBBDDDDDFFFFF1133355577999BBBFBBD5),
    .INIT_17(256'h0000000000000000000000000000B33B5375795557333333111FFFFFFDDDD999),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_008192_004 (
    .addra({addra[10:0],2'b11}),
    .clka(clka),
    .csa(addra[13:11]),
    .dia({open_n1078,open_n1079,open_n1080,open_n1081,open_n1082,4'b0000}),
    .rsta(rsta),
    .doa({open_n1097,open_n1098,open_n1099,open_n1100,open_n1101,inst_doa_i4_007,inst_doa_i4_006,inst_doa_i4_005,inst_doa_i4_004}));
  // address_offset=8192;data_offset=8;depth=1508;width=4;num_section=1;width_per_section=4;section_size=16;working_depth=2048;working_width=4;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("4"),
    .DATA_WIDTH_B("4"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h888881111890333333A11911AAA999222222999933CFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h999A33BFFFFFFFFFFFFFFFFFFFFFF777FFFFFFFF4B9880000008888888888888),
    .INIT_02(256'hFFFFF49000000000888888888888888888089113333111111191AAAA99222A99),
    .INIT_03(256'h800299111111111AAAAA99222199999B33B37FFFFFFFFFFFFFFFFFFF7777FFFF),
    .INIT_04(256'h37FFFFFFFFFFFFFFFFF77777FFFFFFFFFF400000000088888888888888888808),
    .INIT_05(256'h8800000008888888888199999999999111111111111AAAAAA922999999933333),
    .INIT_06(256'h111111AAAAAAAAA19999991333333FFFFFFFFFFFFFFFFFF77777FFFFFFFFFF7F),
    .INIT_07(256'hFFFFFFFFFF777777FFFFFFFF77777E8000000888808808119999999999991111),
    .INIT_08(256'h0888888801111999999999999111111111AAAAAAD6DB99999993333B667FFFFF),
    .INIT_09(256'hAA9EE556591999133356666FFFFFFFFFFFFFFF777777FFFFFFF777777FFE0800),
    .INIT_0A(256'hF7777777FFFF7777777777777708808888891111119999999999991111111AAA),
    .INIT_0B(256'h1111119999999199999111191A1AAD5665665519993BB6E66666FFFFFFFFFFFF),
    .INIT_0C(256'h55E119BBE66666666FFFFFFFFFFF77777777FFF7777777777777777E90888811),
    .INIT_0D(256'hFF77777777777777777FFF088111111111119999999999991111A21D5D555555),
    .INIT_0E(256'h9999999999999911AB6555555555555DA1CE6666666666FFFFFFFFFF77777777),
    .INIT_0F(256'h66666666666FFFFFFFF7777777F77777777777777777777777FE919911111119),
    .INIT_10(256'h77777777EEEEEEEE6E6661111111919999999999991AED65555555555555656E),
    .INIT_11(256'h11A34CC5DD6666666666666666666666666666667FFFFFF77777777777777777),
    .INIT_12(256'h666667FFFF777777777777777777FFEEEEEEEEEEEEEEEEEEE6EE669190819999),
    .INIT_13(256'hEEEEEEEEEEEEE666EEEE6E64BC445DDDDD55DDD5556EEEEE6666666666666666),
    .INIT_14(256'hEE666666666E6EEEEEF77E6666666666667FFF77F7777777777F6EEEEEEEEEEE),
    .INIT_15(256'hF77777777EEEEEEEEEEEEEEEEEEEEEE66EEE666D5DDDDDD55DDDD55DDDD5666E),
    .INIT_16(256'h6E66E6666EEEEE666E6E6666666666666EEEEEEEEE677777FFFFFF77777E666F),
    .INIT_17(256'h00000000000000000000000000007776EEEEE6FFFFF7777777766EEEEEEEEE66),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_008192_008 (
    .addra({addra[10:0],2'b11}),
    .clka(clka),
    .csa(addra[13:11]),
    .dia({open_n1130,open_n1131,open_n1132,open_n1133,open_n1134,4'b0000}),
    .rsta(rsta),
    .doa({open_n1149,open_n1150,open_n1151,open_n1152,open_n1153,inst_doa_i4_011,inst_doa_i4_010,inst_doa_i4_009,inst_doa_i4_008}));
  // address_offset=8192;data_offset=12;depth=1508;width=4;num_section=1;width_per_section=4;section_size=16;working_depth=2048;working_width=4;address_step=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("4"),
    .DATA_WIDTH_B("4"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h555558999667DDDDDDA99999BBB999CCCCCCBBBBEECFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hBBBBEEDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBA6667777775555555555555),
    .INIT_02(256'hFFFFFB677777777755555555555555555556896DDDD999999999BBBB99CCCBBB),
    .INIT_03(256'h567A98999999999BBBBBA9CCCBBBBBBEEEEEFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC77777777755555555555555555565),
    .INIT_05(256'h6677777775555555555766666666669999999999999BBBBBB9CCBBBBBBBEEEEE),
    .INIT_06(256'h999999BBBBBBBBACBBBBBBBEEEEEDEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFEEEEEF6777777555555555886666666666999999),
    .INIT_08(256'h7655555568888666666667999999999999BBBBBBDCBABBBBBBBEEEEBDDFFFFFF),
    .INIT_09(256'hBB9BBCCCEBCBBBBEEEFDDDDEFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEF6677),
    .INIT_0A(256'hFFFFFFFFFFFFFEEEEEEEEEEEEF77675555578888886666666999999999999BBB),
    .INIT_0B(256'h8888887666666A99999999999BCBBCCCCCCCCCCBBBEEEFDDDDDDEFFFFFFFFFFF),
    .INIT_0C(256'hCCBACBDEDEDDDDDDDEFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEF77755588),
    .INIT_0D(256'hFEEEEEEEEEEEEEEEEEEEEF655888888888886666899999999999BCBDCCCCCCCC),
    .INIT_0E(256'h766699999999989ABBCCCCCCCCCCCCCCABEDDDDDDDDDDDEFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hDDDDDDDDDDDEFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEEEEEEEEDD788888888888),
    .INIT_10(256'hEEEEEEEEDCCCCCCCDCDDE7888888876699999999999BCCCCCCCCCCCCCCCCCEDD),
    .INIT_11(256'hA989BAAAAACDDDDDDDDDDDDDDDDDDDDDDDDDDDDDEFFFFFFFFFFFFEEEEEEEEEEE),
    .INIT_12(256'hDDDDDEFFFFFFFFFEEEEEEEEEEEEEEECCCCCCCCCCCCCCCCCCCDCCDE6888699999),
    .INIT_13(256'hCCCCCCCCCCCCCDDDCCCCDCEBABBBBAAAAABBBBBCCCCCCCCCDDDDDDDDDDDDDDDD),
    .INIT_14(256'hCCDDDDDDDDDDDDDDDDDEEDDDDDDDDDDDDDFFFFFFFEEEEEEEEEEEDCCCCCCCCCCC),
    .INIT_15(256'hFFFEEEEEEDCCCCCCCCCCCCCCCCCCCCCDDCCCCCCCCBBBBBBBBBAABBBBBBBCCCCC),
    .INIT_16(256'hDCDDDDDDDCCCCCDDDCDCDDDDDDDDDDDDDDDDDDDDDDEEEEEEEEEEEEFFFFFDDDDE),
    .INIT_17(256'h0000000000000000000000000000FEEDCCCCCDEEEEEEEEEEEEEEEDDDDDDDDDDD),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_9700x16_sub_008192_012 (
    .addra({addra[10:0],2'b11}),
    .clka(clka),
    .csa(addra[13:11]),
    .dia({open_n1182,open_n1183,open_n1184,open_n1185,open_n1186,4'b0000}),
    .rsta(rsta),
    .doa({open_n1201,open_n1202,open_n1203,open_n1204,open_n1205,inst_doa_i4_015,inst_doa_i4_014,inst_doa_i4_013,inst_doa_i4_012}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i0_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i0_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_2  (
    .i0(inst_doa_i4_000),
    .i1(inst_doa_i4_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_3  (
    .i0(inst_doa_i4_000),
    .i1(inst_doa_i4_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b0/B0_2 ),
    .i1(\inst_doa_mux_b0/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b0/B1_0 ),
    .i1(\inst_doa_mux_b0/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i0_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i0_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_2  (
    .i0(inst_doa_i4_001),
    .i1(inst_doa_i4_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_3  (
    .i0(inst_doa_i4_001),
    .i1(inst_doa_i4_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b1/B0_2 ),
    .i1(\inst_doa_mux_b1/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b1/B1_0 ),
    .i1(\inst_doa_mux_b1/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_0  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i0_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_1  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i0_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_2  (
    .i0(inst_doa_i4_010),
    .i1(inst_doa_i4_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_2 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_3  (
    .i0(inst_doa_i4_010),
    .i1(inst_doa_i4_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_3 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b10/B0_0 ),
    .i1(\inst_doa_mux_b10/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b10/B1_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b10/B0_2 ),
    .i1(\inst_doa_mux_b10/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b10/B1_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b10/B1_0 ),
    .i1(\inst_doa_mux_b10/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[10]));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_0  (
    .i0(inst_doa_i0_011),
    .i1(inst_doa_i0_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_1  (
    .i0(inst_doa_i0_011),
    .i1(inst_doa_i0_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_2  (
    .i0(inst_doa_i4_011),
    .i1(inst_doa_i4_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_2 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_3  (
    .i0(inst_doa_i4_011),
    .i1(inst_doa_i4_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_3 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b11/B0_0 ),
    .i1(\inst_doa_mux_b11/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b11/B1_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b11/B0_2 ),
    .i1(\inst_doa_mux_b11/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b11/B1_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b11/B1_0 ),
    .i1(\inst_doa_mux_b11/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[11]));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_0  (
    .i0(inst_doa_i0_012),
    .i1(inst_doa_i0_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_0 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_1  (
    .i0(inst_doa_i0_012),
    .i1(inst_doa_i0_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_1 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_2  (
    .i0(inst_doa_i4_012),
    .i1(inst_doa_i4_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_2 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_3  (
    .i0(inst_doa_i4_012),
    .i1(inst_doa_i4_012),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_3 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b12/B0_0 ),
    .i1(\inst_doa_mux_b12/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b12/B1_0 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b12/B0_2 ),
    .i1(\inst_doa_mux_b12/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b12/B1_1 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b12/B1_0 ),
    .i1(\inst_doa_mux_b12/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[12]));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_0  (
    .i0(inst_doa_i0_013),
    .i1(inst_doa_i0_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_0 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_1  (
    .i0(inst_doa_i0_013),
    .i1(inst_doa_i0_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_1 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_2  (
    .i0(inst_doa_i4_013),
    .i1(inst_doa_i4_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_2 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_3  (
    .i0(inst_doa_i4_013),
    .i1(inst_doa_i4_013),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_3 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b13/B0_0 ),
    .i1(\inst_doa_mux_b13/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b13/B1_0 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b13/B0_2 ),
    .i1(\inst_doa_mux_b13/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b13/B1_1 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b13/B1_0 ),
    .i1(\inst_doa_mux_b13/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[13]));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_0  (
    .i0(inst_doa_i0_014),
    .i1(inst_doa_i0_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_0 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_1  (
    .i0(inst_doa_i0_014),
    .i1(inst_doa_i0_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_1 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_2  (
    .i0(inst_doa_i4_014),
    .i1(inst_doa_i4_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_2 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_3  (
    .i0(inst_doa_i4_014),
    .i1(inst_doa_i4_014),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_3 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b14/B0_0 ),
    .i1(\inst_doa_mux_b14/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b14/B1_0 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b14/B0_2 ),
    .i1(\inst_doa_mux_b14/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b14/B1_1 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b14/B1_0 ),
    .i1(\inst_doa_mux_b14/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[14]));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_0  (
    .i0(inst_doa_i0_015),
    .i1(inst_doa_i0_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_0 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_1  (
    .i0(inst_doa_i0_015),
    .i1(inst_doa_i0_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_1 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_2  (
    .i0(inst_doa_i4_015),
    .i1(inst_doa_i4_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_2 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_3  (
    .i0(inst_doa_i4_015),
    .i1(inst_doa_i4_015),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_3 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b15/B0_0 ),
    .i1(\inst_doa_mux_b15/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b15/B1_0 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b15/B0_2 ),
    .i1(\inst_doa_mux_b15/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b15/B1_1 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b15/B1_0 ),
    .i1(\inst_doa_mux_b15/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[15]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i0_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i0_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_2  (
    .i0(inst_doa_i4_002),
    .i1(inst_doa_i4_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_3  (
    .i0(inst_doa_i4_002),
    .i1(inst_doa_i4_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b2/B0_2 ),
    .i1(\inst_doa_mux_b2/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b2/B1_0 ),
    .i1(\inst_doa_mux_b2/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i0_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i0_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_2  (
    .i0(inst_doa_i4_003),
    .i1(inst_doa_i4_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_2 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_3  (
    .i0(inst_doa_i4_003),
    .i1(inst_doa_i4_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_3 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b3/B0_2 ),
    .i1(\inst_doa_mux_b3/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b3/B1_0 ),
    .i1(\inst_doa_mux_b3/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i0_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i0_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_2  (
    .i0(inst_doa_i4_004),
    .i1(inst_doa_i4_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_2 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_3  (
    .i0(inst_doa_i4_004),
    .i1(inst_doa_i4_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_3 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b4/B0_2 ),
    .i1(\inst_doa_mux_b4/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b4/B1_0 ),
    .i1(\inst_doa_mux_b4/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i0_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i0_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_2  (
    .i0(inst_doa_i4_005),
    .i1(inst_doa_i4_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_2 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_3  (
    .i0(inst_doa_i4_005),
    .i1(inst_doa_i4_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_3 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b5/B0_2 ),
    .i1(\inst_doa_mux_b5/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b5/B1_0 ),
    .i1(\inst_doa_mux_b5/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i0_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i0_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_2  (
    .i0(inst_doa_i4_006),
    .i1(inst_doa_i4_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_2 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_3  (
    .i0(inst_doa_i4_006),
    .i1(inst_doa_i4_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_3 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b6/B0_2 ),
    .i1(\inst_doa_mux_b6/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b6/B1_0 ),
    .i1(\inst_doa_mux_b6/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i0_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i0_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_2  (
    .i0(inst_doa_i4_007),
    .i1(inst_doa_i4_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_2 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_3  (
    .i0(inst_doa_i4_007),
    .i1(inst_doa_i4_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_3 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b7/B0_2 ),
    .i1(\inst_doa_mux_b7/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b7/B1_0 ),
    .i1(\inst_doa_mux_b7/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[7]));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_0  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i0_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_1  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i0_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_2  (
    .i0(inst_doa_i4_008),
    .i1(inst_doa_i4_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_2 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_3  (
    .i0(inst_doa_i4_008),
    .i1(inst_doa_i4_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_3 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b8/B0_0 ),
    .i1(\inst_doa_mux_b8/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b8/B0_2 ),
    .i1(\inst_doa_mux_b8/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b8/B1_0 ),
    .i1(\inst_doa_mux_b8/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[8]));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_0  (
    .i0(inst_doa_i0_009),
    .i1(inst_doa_i0_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_1  (
    .i0(inst_doa_i0_009),
    .i1(inst_doa_i0_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_2  (
    .i0(inst_doa_i4_009),
    .i1(inst_doa_i4_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_2 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_3  (
    .i0(inst_doa_i4_009),
    .i1(inst_doa_i4_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_3 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b9/B0_0 ),
    .i1(\inst_doa_mux_b9/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b9/B1_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b9/B0_2 ),
    .i1(\inst_doa_mux_b9/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b9/B1_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b9/B1_0 ),
    .i1(\inst_doa_mux_b9/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[9]));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

